`define ALU_1   'h8
`define ALU_2   'h9
`define ALU_ADD 'hA
`define ALU_SUB 'hB
`define ALU_RS  'hC
`define ALU_LS  'hD
`define ALU_AND 'hE
`define ALU_OR  'hF
`define ALU_NOT 'h10
`define ALU_GT  'h11
`define ALU_LT  'h12
`define ALU_EQ  'h13
`define ALU_OV  'h14

`define IO_INP1 'h1000
`define IO_INP2 'h1001
`define IO_INP3 'h1002
`define IO_OUT1 'h1003
`define IO_OUT2 'h1004
`define IO_OUT3 'h1005
`define IO_POP  'h1006

`define VRAM_START 'h1800
`define VRAM_END   'h1C00

`define RAM_START 'h4000
`define RAM_END   'hFFFF
