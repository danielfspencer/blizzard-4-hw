`define WORD_SIZE 16
`define WORD [`WORD_SIZE - 1:0]
