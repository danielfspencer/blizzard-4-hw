`define CLOCKS input reset, \
    input read_clk, \
    input write_clk, \
    input ctrl_clk
